correct_real[0] = 32'sd0; correct_imag[0] = 32'h0;
correct_real[1] = 32'sd70; correct_imag[1] = -32'h1434;
correct_real[2] = 32'sd281; correct_imag[2] = -32'h2856;
correct_real[3] = 32'sd659; correct_imag[3] = -32'h4445;
correct_real[4] = 32'sd1286; correct_imag[4] = -32'h6465;
correct_real[5] = 32'sd5831; correct_imag[5] = -32'h23281;
correct_real[6] = 32'sd2113; correct_imag[6] = -32'h6968;
correct_real[7] = 32'sd3399; correct_imag[7] = -32'h9501;
correct_real[8] = 32'sd4862; correct_imag[8] = -32'h11738;
correct_real[9] = 32'sd6691; correct_imag[9] = -32'h14148;
correct_real[10] = 32'sd9033; correct_imag[10] = -32'h16900;
correct_real[11] = 32'sd12119; correct_imag[11] = -32'h20219;
correct_real[12] = 32'sd16293; correct_imag[12] = -32'h24384;
correct_real[13] = 32'sd22166; correct_imag[13] = -32'h29888;
correct_real[14] = 32'sd30930; correct_imag[14] = -32'h37688;
correct_real[15] = 32'sd45234; correct_imag[15] = -32'h49908;
correct_real[16] = 32'sd72330; correct_imag[16] = -32'h72330;
correct_real[17] = 32'sd142090; correct_imag[17] = -32'h128783;
correct_real[18] = 32'sd702518; correct_imag[18] = -32'h576542;
correct_real[19] = -32'sd307234; correct_imag[19] = 32'h227860;
correct_real[20] = -32'sd139371; correct_imag[20] = 32'h93125;
correct_real[21] = -32'sd95491; correct_imag[21] = 32'h57235;
correct_real[22] = -32'sd75464; correct_imag[22] = 32'h40336;
correct_real[23] = -32'sd64138; correct_imag[23] = 32'h30335;
correct_real[24] = -32'sd56956; correct_imag[24] = 32'h23591;
correct_real[25] = -32'sd52082; correct_imag[25] = 32'h18635;
correct_real[26] = -32'sd48648; correct_imag[26] = 32'h14757;
correct_real[27] = -32'sd46168; correct_imag[27] = 32'h11564;
correct_real[28] = -32'sd44379; correct_imag[28] = 32'h8827;
correct_real[29] = -32'sd43109; correct_imag[29] = 32'h6394;
correct_real[30] = -32'sd42268; correct_imag[30] = 32'h4163;
correct_real[31] = -32'sd41783; correct_imag[31] = 32'h2052;
correct_real[32] = -32'sd41632; correct_imag[32] = 32'h0;
correct_real[33] = -32'sd41783; correct_imag[33] = -32'h2052;
correct_real[34] = -32'sd42268; correct_imag[34] = -32'h4163;
correct_real[35] = -32'sd43109; correct_imag[35] = -32'h6394;
correct_real[36] = -32'sd44379; correct_imag[36] = -32'h8827;
correct_real[37] = -32'sd46168; correct_imag[37] = -32'h11564;
correct_real[38] = -32'sd48648; correct_imag[38] = -32'h14757;
correct_real[39] = -32'sd52082; correct_imag[39] = -32'h18635;
correct_real[40] = -32'sd56956; correct_imag[40] = -32'h23591;
correct_real[41] = -32'sd64138; correct_imag[41] = -32'h30335;
correct_real[42] = -32'sd75464; correct_imag[42] = -32'h40336;
correct_real[43] = -32'sd95491; correct_imag[43] = -32'h57235;
correct_real[44] = -32'sd139371; correct_imag[44] = -32'h93125;
correct_real[45] = -32'sd307234; correct_imag[45] = -32'h227860;
correct_real[46] = 32'sd702518; correct_imag[46] = 32'h576542;
correct_real[47] = 32'sd142090; correct_imag[47] = 32'h128783;
correct_real[48] = 32'sd72330; correct_imag[48] = 32'h72330;
correct_real[49] = 32'sd45234; correct_imag[49] = 32'h49908;
correct_real[50] = 32'sd30930; correct_imag[50] = 32'h37688;
correct_real[51] = 32'sd22166; correct_imag[51] = 32'h29888;
correct_real[52] = 32'sd16293; correct_imag[52] = 32'h24384;
correct_real[53] = 32'sd12119; correct_imag[53] = 32'h20219;
correct_real[54] = 32'sd9033; correct_imag[54] = 32'h16900;
correct_real[55] = 32'sd6691; correct_imag[55] = 32'h14148;
correct_real[56] = 32'sd4862; correct_imag[56] = 32'h11738;
correct_real[57] = 32'sd3399; correct_imag[57] = 32'h9501;
correct_real[58] = 32'sd2113; correct_imag[58] = 32'h6968;
correct_real[59] = 32'sd5831; correct_imag[59] = 32'h23281;
correct_real[60] = 32'sd1286; correct_imag[60] = 32'h6465;
correct_real[61] = 32'sd659; correct_imag[61] = 32'h4445;
correct_real[62] = 32'sd281; correct_imag[62] = 32'h2856;
correct_real[63] = 32'sd70; correct_imag[63] = 32'h1434;
