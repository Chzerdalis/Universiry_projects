w_real[0] = 16'h7FFF; w_imag[0] = 16'h0000;
w_real[1] = 16'h7F62; w_imag[1] = 16'hF375;
w_real[2] = 16'h7D8A; w_imag[2] = 16'hE708;
w_real[3] = 16'h7A7D; w_imag[3] = 16'hDAD8;
w_real[4] = 16'h7641; w_imag[4] = 16'hCF05;
w_real[5] = 16'h70E2; w_imag[5] = 16'hC3AA;
w_real[6] = 16'h6A6D; w_imag[6] = 16'hB8E4;
w_real[7] = 16'h62F2; w_imag[7] = 16'hAECD;
w_real[8] = 16'h5A82; w_imag[8] = 16'hA57E;
w_real[9] = 16'h5133; w_imag[9] = 16'h9D0E;
w_real[10] = 16'h471C; w_imag[10] = 16'h9593;
w_real[11] = 16'h3C56; w_imag[11] = 16'h8F1E;
w_real[12] = 16'h30FB; w_imag[12] = 16'h89BF;
w_real[13] = 16'h2528; w_imag[13] = 16'h8583;
w_real[14] = 16'h18F8; w_imag[14] = 16'h8276;
w_real[15] = 16'h0C8B; w_imag[15] = 16'h809E;
w_real[16] = 16'h0000; w_imag[16] = 16'h8000;
w_real[17] = 16'hF375; w_imag[17] = 16'h809E;
w_real[18] = 16'hE708; w_imag[18] = 16'h8276;
w_real[19] = 16'hDAD8; w_imag[19] = 16'h8583;
w_real[20] = 16'hCF05; w_imag[20] = 16'h89BF;
w_real[21] = 16'hC3AA; w_imag[21] = 16'h8F1E;
w_real[22] = 16'hB8E4; w_imag[22] = 16'h9593;
w_real[23] = 16'hAECD; w_imag[23] = 16'h9D0E;
w_real[24] = 16'hA57E; w_imag[24] = 16'hA57E;
w_real[25] = 16'h9D0E; w_imag[25] = 16'hAECD;
w_real[26] = 16'h9593; w_imag[26] = 16'hB8E4;
w_real[27] = 16'h8F1E; w_imag[27] = 16'hC3AA;
w_real[28] = 16'h89BF; w_imag[28] = 16'hCF05;
w_real[29] = 16'h8583; w_imag[29] = 16'hDAD8;
w_real[30] = 16'h8276; w_imag[30] = 16'hE708;
w_real[31] = 16'h809E; w_imag[31] = 16'hF375;
w_real[32] = 16'h8000; w_imag[32] = 16'h0000;
w_real[33] = 16'h809E; w_imag[33] = 16'h0C8B;
w_real[34] = 16'h8276; w_imag[34] = 16'h18F8;
w_real[35] = 16'h8583; w_imag[35] = 16'h2528;
w_real[36] = 16'h89BF; w_imag[36] = 16'h30FB;
w_real[37] = 16'h8F1E; w_imag[37] = 16'h3C56;
w_real[38] = 16'h9593; w_imag[38] = 16'h471C;
w_real[39] = 16'h9D0E; w_imag[39] = 16'h5133;
w_real[40] = 16'hA57E; w_imag[40] = 16'h5A82;
w_real[41] = 16'hAECD; w_imag[41] = 16'h62F2;
w_real[42] = 16'hB8E4; w_imag[42] = 16'h6A6D;
w_real[43] = 16'hC3AA; w_imag[43] = 16'h70E2;
w_real[44] = 16'hCF05; w_imag[44] = 16'h7641;
w_real[45] = 16'hDAD8; w_imag[45] = 16'h7A7D;
w_real[46] = 16'hE708; w_imag[46] = 16'h7D8A;
w_real[47] = 16'hF375; w_imag[47] = 16'h7F62;
w_real[48] = 16'h0000; w_imag[48] = 16'h7FFF;
w_real[49] = 16'h0C8B; w_imag[49] = 16'h7F62;
w_real[50] = 16'h18F8; w_imag[50] = 16'h7D8A;
w_real[51] = 16'h2528; w_imag[51] = 16'h7A7D;
w_real[52] = 16'h30FB; w_imag[52] = 16'h7641;
w_real[53] = 16'h3C56; w_imag[53] = 16'h70E2;
w_real[54] = 16'h471C; w_imag[54] = 16'h6A6D;
w_real[55] = 16'h5133; w_imag[55] = 16'h62F2;
w_real[56] = 16'h5A82; w_imag[56] = 16'h5A82;
w_real[57] = 16'h62F2; w_imag[57] = 16'h5133;
w_real[58] = 16'h6A6D; w_imag[58] = 16'h471C;
w_real[59] = 16'h70E2; w_imag[59] = 16'h3C56;
w_real[60] = 16'h7641; w_imag[60] = 16'h30FB;
w_real[61] = 16'h7A7D; w_imag[61] = 16'h2528;
w_real[62] = 16'h7D8A; w_imag[62] = 16'h18F8;
w_real[63] = 16'h7F62; w_imag[63] = 16'h0C8B;
