input_real_arr[0] = 32'sd0;
input_real_arr[32] = 32'sd32767;
input_real_arr[16] = -32'sd6738;
input_real_arr[48] = -32'sd24327;
input_real_arr[8] = 32'sd9756;
input_real_arr[40] = 32'sd15217;
input_real_arr[24] = -32'sd10062;
input_real_arr[56] = -32'sd7920;
input_real_arr[4] = 32'sd10717;
input_real_arr[36] = 32'sd3571;
input_real_arr[20] = -32'sd11792;
input_real_arr[52] = -32'sd1924;
input_real_arr[12] = 32'sd10901;
input_real_arr[44] = 32'sd958;
input_real_arr[28] = -32'sd7267;
input_real_arr[60] = -32'sd1439;
input_real_arr[2] = 32'sd2208;
input_real_arr[34] = 32'sd2554;
input_real_arr[18] = 32'sd2413;
input_real_arr[50] = -32'sd1936;
input_real_arr[10] = -32'sd4438;
input_real_arr[42] = -32'sd699;
input_real_arr[26] = 32'sd4139;
input_real_arr[58] = 32'sd4303;
input_real_arr[6] = -32'sd3791;
input_real_arr[38] = -32'sd6510;
input_real_arr[22] = 32'sd3481;
input_real_arr[54] = 32'sd4526;
input_real_arr[14] = -32'sd2133;
input_real_arr[46] = 32'sd594;
input_real_arr[30] = -32'sd783;
input_real_arr[62] = -32'sd3037;
input_real_arr[1] = 32'sd3037;
input_real_arr[33] = 32'sd783;
input_real_arr[17] = -32'sd594;
input_real_arr[49] = 32'sd2133;
input_real_arr[9] = -32'sd4526;
input_real_arr[41] = -32'sd3481;
input_real_arr[25] = 32'sd6510;
input_real_arr[57] = 32'sd3791;
input_real_arr[5] = -32'sd4303;
input_real_arr[37] = -32'sd4139;
input_real_arr[21] = 32'sd699;
input_real_arr[53] = 32'sd4438;
input_real_arr[13] = 32'sd1936;
input_real_arr[45] = -32'sd2413;
input_real_arr[29] = -32'sd2554;
input_real_arr[61] = -32'sd2208;
input_real_arr[3] = 32'sd1439;
input_real_arr[35] = 32'sd7267;
input_real_arr[19] = -32'sd958;
input_real_arr[51] = -32'sd10901;
input_real_arr[11] = 32'sd1924;
input_real_arr[43] = 32'sd11792;
input_real_arr[27] = -32'sd3571;
input_real_arr[59] = -32'sd10717;
input_real_arr[7] = 32'sd7920;
input_real_arr[39] = 32'sd10062;
input_real_arr[23] = -32'sd15217;
input_real_arr[55] = -32'sd9756;
input_real_arr[15] = 32'sd24327;
input_real_arr[47] = 32'sd6738;
input_real_arr[31] = -32'sd32767;
input_real_arr[63] = 32'sd0;
