`timescale 1ns/1ps

module vram_red(reset, clk, address, red);
    input clk, reset;
    input [13:0] address;
    output red;
    wire input_data, ram_enable, reg_enable, write_enable;

    assign input_data = 0;
    assign ram_enable = 1'b1;
    assign reg_enable = 0;
    assign write_enable = 0;

    BRAM_SINGLE_MACRO #(
        .BRAM_SIZE("18Kb"), // Target BRAM, "18Kb" or "36Kb" 
        .DEVICE("7SERIES"), // Target Device: "7SERIES" 
        .DO_REG(0), // Optional output register (0 or 1)
        .INIT(36'h000000000), // Initial values on output port
        .INIT_FILE ("NONE"),
        .WRITE_WIDTH(1), // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        .READ_WIDTH(1),  // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        .SRVAL(36'h000000000), // Set/Reset value for port output
        .WRITE_MODE("READ_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
        
        .INIT_00(256'hffffffffffffffffffffffffffffffff_ffffffffffffffffffffffffffffffff),
        .INIT_01(256'hffffffffffffffffffffffffffffffff_ffffffffffffffffffffffffffffffff),
        .INIT_02(256'hffffffffffffffffffffffffffffffff_ffffffffffffffffffffffffffffffff),
        .INIT_03(256'hffffffffffffffffffffffffffffffff_ffffffffffffffffffffffffffffffff),
        .INIT_04(256'hffffc7fffffffff01fffffffffffffff_ffff00003fffffc007ffffffffffffff),
        .INIT_05(256'hfffe00001fffff8003ffffffffffffff_fffe00000fffff0001ffffffffffffff),
        .INIT_06(256'hfffe000007fffe0000ffffffffffffff_fffe000003fffc00007fffffffffffff),
        .INIT_07(256'hfffe000007fffc00007fffffffffffff_fffe00000ffff800003fffffffffffff),
        .INIT_08(256'hfffe000007fff800003fffffffffffff_fffe000007fff800003fffffffffffff),
        .INIT_09(256'hfffe000003fff800003fffffffffffff_fffe000003fff800003fffffffffffff),
        .INIT_0A(256'hfffe000003fff800003fffffffffffff_fffe000003fff800003fffffffffffff),
        .INIT_0B(256'hfffe000003fffc00007fffffffffffff_fffe000003fffc00007fffffffffffff),
        .INIT_0C(256'hfffe000003fffe0000ffffffffffffff_fffe000003ffff0001ffffffffffffff),
        .INIT_0D(256'hfffe000003ffff8003ffffffffffffff_fffe000003ffffc007ffffffffffffff),
        .INIT_0E(256'hfffe000003fffff01fffffffffffffff_fffe000003fffffc7fffffffffffffff),
        .INIT_0F(256'hfffe000003fffffc7fffffffffffffff_fffe000003fffffc7fffffffffffffff),
        .INIT_10(256'hfffe000003fffffc7fffffffffffffff_fffe000007fffffc7fffffffffffffff),
        .INIT_11(256'hffff07fffffffffc7fffffffffffffff_fffffffffffffffc7fffffffffffffff),
        .INIT_12(256'hfffffffffffffffc7fffffffffffffff_fffffffffffffffc7fffffffffffffff),
        .INIT_13(256'hfffffffffffffffc7fffffffffffffff_fffffffffffffffc7fffffffffffffff),
        .INIT_14(256'hfffffffffffffffc7fffffffffffffff_fffffffffffffffc7fffffffffffffff),
        .INIT_15(256'hfffffffffffffffc7fffffffffffffff_fffffffffffffffc7fffffffffffffff),
        .INIT_16(256'hfffffffffffffffc7fffffffffffffff_fffffffffffffffc7fffffffffffffff),
        .INIT_17(256'hfffffffffffffffc7fffffffffffffff_fffffffffffffffc7fffffffffffffff),
        .INIT_18(256'hfffffffffffffff83fffffffffffffff_fffffffffffffff81fffffffffffffff),
        .INIT_19(256'hfffffffffffffff00fffffffffffffff_ffffffffffffffe007ffffffffffffff),
        .INIT_1A(256'hffffffffffffff8003ffffffffffffff_ffffffffffffff0441ffffffffffffff),
        .INIT_1B(256'hfffffffffffffe0c60ffffffffffffff_fffffffffffffc1c707fffffffffffff),
        .INIT_1C(256'hfffffffffffff83c783fffffffffffff_fffffffffffff07c7c1fffffffffffff),
        .INIT_1D(256'hffffffffffffe0fc7e0fffffffffffff_ffffffffffffc1fc7f07ffffffffffff),
        .INIT_1E(256'hffffffffffff83fc7f83ffffffffffff_ffffffffffff07fc7fc1ffffffffffff),
        .INIT_1F(256'hfffffffffffe0ffc7fe0ffffffffffff_fffffffffffc1ffc7ff07fffffffffff),
        .INIT_20(256'hfffffffffff83ffc7ff83fffffffffff_fffffffffff07ffc7ffc1fffffffffff),
        .INIT_21(256'hffffffffffe0fffc7ffe0fffffffffff_ffffffffffc1fffc7fff07ffffffffff),
        .INIT_22(256'hffffffffffe3fffc7fff8fffffffffff_fffffffffff7fffc7fffdfffffffffff),
        .INIT_23(256'hfffffffffffffffc7fffffffffffffff_fffffffffffffffc7fffffffffffffff),
        .INIT_24(256'hfffffffffffffffc7fffffffffffffff_fffffffffffffffc7fffffffffffffff),
        .INIT_25(256'hfffffffffffffffc7fffffffffffffff_fffffffffffffffc7fffffffffffffff),
        .INIT_26(256'hfffffffffffffffc7fffffffffffffff_fffffffffffffffc7fffffffffffffff),
        .INIT_27(256'hfffffffffffffff83fffffffffffffff_fffffffffffffff01fffffffffffffff),
        .INIT_28(256'hffffffffffffffe00fffffffffffffff_ffffffffffffffc107ffffffffffffff),
        .INIT_29(256'hffffffffffffff8383ffffffffffffff_ffffffffffffff07c1ffffffffffffff),
        .INIT_2A(256'hfffffffffffffe0fe0ffffffffffffff_fffffffffffffc1ff07fffffffffffff),
        .INIT_2B(256'hfffffffffffff83ff83fffffffffffff_fffffffffffff07ffc1fffffffffffff),
        .INIT_2C(256'hffffffffffffe0fffe0fffffffffffff_ffffffffffffc1ffff07ffffffffffff),
        .INIT_2D(256'hffffffffffff83ffff83ffffffffffff_ffffffffffff07ffffc1ffffffffffff),
        .INIT_2E(256'hfffffffffffe0fffffe0ffffffffffff_fffffffffffc1ffffff07fffffffffff),
        .INIT_2F(256'hfffffffffff83ffffff83fffffffffff_fffffffffff07ffffffc1fffffffffff)   
    ) BRAM_SINGLE_MACRO_inst (
        .DO(red),       // Output data, width defined by READ_WIDTH parameter
        .ADDR(address),   // Input address, width defined by read/write port depth
        .CLK(clk),     // 1-bit input clock
        .DI(input_data),       // Input data port, width defined by WRITE_WIDTH parameter
        .EN(ram_enable),       // 1-bit input RAM enable
        .REGCE(reg_enable), // 1-bit input output register enable
        .RST(reset),     // 1-bit input reset
        .WE(write_enable)        // Input write enable, width defined by write port depth
    );								
endmodule