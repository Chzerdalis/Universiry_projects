input_real_arr[0] = 32'sd0;
input_real_arr[128] = 32'sd32767;
input_real_arr[64] = -32'sd609;
input_real_arr[192] = -32'sd26021;
input_real_arr[32] = 32'sd1595;
input_real_arr[160] = 32'sd19510;
input_real_arr[96] = -32'sd2729;
input_real_arr[224] = -32'sd15929;
input_real_arr[16] = 32'sd3910;
input_real_arr[144] = 32'sd13024;
input_real_arr[80] = -32'sd5655;
input_real_arr[208] = -32'sd9141;
input_real_arr[48] = 32'sd7846;
input_real_arr[176] = 32'sd6167;
input_real_arr[112] = -32'sd9500;
input_real_arr[240] = -32'sd7089;
input_real_arr[8] = 32'sd9488;
input_real_arr[136] = 32'sd10326;
input_real_arr[72] = -32'sd8186;
input_real_arr[200] = -32'sd11345;
input_real_arr[40] = 32'sd7997;
input_real_arr[168] = 32'sd7976;
input_real_arr[104] = -32'sd9273;
input_real_arr[232] = -32'sd1727;
input_real_arr[24] = 32'sd9925;
input_real_arr[152] = -32'sd3975;
input_real_arr[88] = -32'sd9835;
input_real_arr[216] = 32'sd8019;
input_real_arr[56] = 32'sd10199;
input_real_arr[184] = -32'sd11693;
input_real_arr[120] = -32'sd11091;
input_real_arr[248] = 32'sd14416;
input_real_arr[4] = 32'sd11988;
input_real_arr[132] = -32'sd13998;
input_real_arr[68] = -32'sd12181;
input_real_arr[196] = 32'sd9912;
input_real_arr[36] = 32'sd11092;
input_real_arr[164] = -32'sd4816;
input_real_arr[100] = -32'sd9045;
input_real_arr[228] = 32'sd1870;
input_real_arr[20] = 32'sd7881;
input_real_arr[148] = -32'sd960;
input_real_arr[84] = -32'sd8876;
input_real_arr[212] = 32'sd981;
input_real_arr[52] = 32'sd10036;
input_real_arr[180] = -32'sd2148;
input_real_arr[116] = -32'sd9601;
input_real_arr[244] = 32'sd4378;
input_real_arr[12] = 32'sd8752;
input_real_arr[140] = -32'sd6791;
input_real_arr[76] = -32'sd8600;
input_real_arr[204] = 32'sd7467;
input_real_arr[44] = 32'sd8475;
input_real_arr[172] = -32'sd5095;
input_real_arr[108] = -32'sd6795;
input_real_arr[236] = 32'sd1691;
input_real_arr[28] = 32'sd3832;
input_real_arr[156] = 32'sd376;
input_real_arr[92] = -32'sd1674;
input_real_arr[220] = -32'sd2009;
input_real_arr[60] = 32'sd653;
input_real_arr[188] = 32'sd4037;
input_real_arr[124] = -32'sd341;
input_real_arr[252] = -32'sd4453;
input_real_arr[2] = 32'sd875;
input_real_arr[130] = 32'sd1931;
input_real_arr[66] = -32'sd1192;
input_real_arr[194] = 32'sd1810;
input_real_arr[34] = 32'sd589;
input_real_arr[162] = -32'sd4431;
input_real_arr[98] = 32'sd374;
input_real_arr[226] = 32'sd5559;
input_real_arr[18] = -32'sd1745;
input_real_arr[146] = -32'sd5947;
input_real_arr[82] = 32'sd3476;
input_real_arr[210] = 32'sd5442;
input_real_arr[50] = -32'sd4925;
input_real_arr[178] = -32'sd3857;
input_real_arr[114] = 32'sd5750;
input_real_arr[242] = 32'sd2133;
input_real_arr[10] = -32'sd5403;
input_real_arr[138] = -32'sd792;
input_real_arr[74] = 32'sd3434;
input_real_arr[202] = -32'sd351;
input_real_arr[42] = -32'sd532;
input_real_arr[170] = 32'sd500;
input_real_arr[106] = -32'sd2004;
input_real_arr[234] = 32'sd1075;
input_real_arr[26] = 32'sd3657;
input_real_arr[154] = -32'sd3291;
input_real_arr[90] = -32'sd4571;
input_real_arr[218] = 32'sd4840;
input_real_arr[58] = 32'sd4339;
input_real_arr[186] = -32'sd5620;
input_real_arr[122] = -32'sd3003;
input_real_arr[250] = 32'sd5607;
input_real_arr[6] = 32'sd2161;
input_real_arr[134] = -32'sd4811;
input_real_arr[70] = -32'sd2944;
input_real_arr[198] = 32'sd4203;
input_real_arr[38] = 32'sd4408;
input_real_arr[166] = -32'sd3927;
input_real_arr[102] = -32'sd5486;
input_real_arr[230] = 32'sd2978;
input_real_arr[22] = 32'sd6757;
input_real_arr[150] = -32'sd2013;
input_real_arr[86] = -32'sd8781;
input_real_arr[214] = 32'sd2948;
input_real_arr[54] = 32'sd9985;
input_real_arr[182] = -32'sd6257;
input_real_arr[118] = -32'sd8370;
input_real_arr[246] = 32'sd10089;
input_real_arr[14] = 32'sd4647;
input_real_arr[142] = -32'sd12025;
input_real_arr[78] = -32'sd728;
input_real_arr[206] = 32'sd12023;
input_real_arr[46] = -32'sd2476;
input_real_arr[174] = -32'sd12135;
input_real_arr[110] = 32'sd4149;
input_real_arr[238] = 32'sd12914;
input_real_arr[30] = -32'sd4742;
input_real_arr[158] = -32'sd12215;
input_real_arr[94] = 32'sd5909;
input_real_arr[222] = 32'sd8806;
input_real_arr[62] = -32'sd6892;
input_real_arr[190] = -32'sd5075;
input_real_arr[126] = 32'sd5852;
input_real_arr[254] = 32'sd4183;
input_real_arr[1] = -32'sd4183;
input_real_arr[129] = -32'sd5852;
input_real_arr[65] = 32'sd5075;
input_real_arr[193] = 32'sd6892;
input_real_arr[33] = -32'sd8806;
input_real_arr[161] = -32'sd5909;
input_real_arr[97] = 32'sd12215;
input_real_arr[225] = 32'sd4742;
input_real_arr[17] = -32'sd12914;
input_real_arr[145] = -32'sd4149;
input_real_arr[81] = 32'sd12135;
input_real_arr[209] = 32'sd2476;
input_real_arr[49] = -32'sd12023;
input_real_arr[177] = 32'sd728;
input_real_arr[113] = 32'sd12025;
input_real_arr[241] = -32'sd4647;
input_real_arr[9] = -32'sd10089;
input_real_arr[137] = 32'sd8370;
input_real_arr[73] = 32'sd6257;
input_real_arr[201] = -32'sd9985;
input_real_arr[41] = -32'sd2948;
input_real_arr[169] = 32'sd8781;
input_real_arr[105] = 32'sd2013;
input_real_arr[233] = -32'sd6757;
input_real_arr[25] = -32'sd2978;
input_real_arr[153] = 32'sd5486;
input_real_arr[89] = 32'sd3927;
input_real_arr[217] = -32'sd4408;
input_real_arr[57] = -32'sd4203;
input_real_arr[185] = 32'sd2944;
input_real_arr[121] = 32'sd4811;
input_real_arr[249] = -32'sd2161;
input_real_arr[5] = -32'sd5607;
input_real_arr[133] = 32'sd3003;
input_real_arr[69] = 32'sd5620;
input_real_arr[197] = -32'sd4339;
input_real_arr[37] = -32'sd4840;
input_real_arr[165] = 32'sd4571;
input_real_arr[101] = 32'sd3291;
input_real_arr[229] = -32'sd3657;
input_real_arr[21] = -32'sd1075;
input_real_arr[149] = 32'sd2004;
input_real_arr[85] = -32'sd500;
input_real_arr[213] = 32'sd532;
input_real_arr[53] = 32'sd351;
input_real_arr[181] = -32'sd3434;
input_real_arr[117] = 32'sd792;
input_real_arr[245] = 32'sd5403;
input_real_arr[13] = -32'sd2133;
input_real_arr[141] = -32'sd5750;
input_real_arr[77] = 32'sd3857;
input_real_arr[205] = 32'sd4925;
input_real_arr[45] = -32'sd5442;
input_real_arr[173] = -32'sd3476;
input_real_arr[109] = 32'sd5947;
input_real_arr[237] = 32'sd1745;
input_real_arr[29] = -32'sd5559;
input_real_arr[157] = -32'sd374;
input_real_arr[93] = 32'sd4431;
input_real_arr[221] = -32'sd589;
input_real_arr[61] = -32'sd1810;
input_real_arr[189] = 32'sd1192;
input_real_arr[125] = -32'sd1931;
input_real_arr[253] = -32'sd875;
input_real_arr[3] = 32'sd4453;
input_real_arr[131] = 32'sd341;
input_real_arr[67] = -32'sd4037;
input_real_arr[195] = -32'sd653;
input_real_arr[35] = 32'sd2009;
input_real_arr[163] = 32'sd1674;
input_real_arr[99] = -32'sd376;
input_real_arr[227] = -32'sd3832;
input_real_arr[19] = -32'sd1691;
input_real_arr[147] = 32'sd6795;
input_real_arr[83] = 32'sd5095;
input_real_arr[211] = -32'sd8475;
input_real_arr[51] = -32'sd7467;
input_real_arr[179] = 32'sd8600;
input_real_arr[115] = 32'sd6791;
input_real_arr[243] = -32'sd8752;
input_real_arr[11] = -32'sd4378;
input_real_arr[139] = 32'sd9601;
input_real_arr[75] = 32'sd2148;
input_real_arr[203] = -32'sd10036;
input_real_arr[43] = -32'sd981;
input_real_arr[171] = 32'sd8876;
input_real_arr[107] = 32'sd960;
input_real_arr[235] = -32'sd7881;
input_real_arr[27] = -32'sd1870;
input_real_arr[155] = 32'sd9045;
input_real_arr[91] = 32'sd4816;
input_real_arr[219] = -32'sd11092;
input_real_arr[59] = -32'sd9912;
input_real_arr[187] = 32'sd12181;
input_real_arr[123] = 32'sd13998;
input_real_arr[251] = -32'sd11988;
input_real_arr[7] = -32'sd14416;
input_real_arr[135] = 32'sd11091;
input_real_arr[71] = 32'sd11693;
input_real_arr[199] = -32'sd10199;
input_real_arr[39] = -32'sd8019;
input_real_arr[167] = 32'sd9835;
input_real_arr[103] = 32'sd3975;
input_real_arr[231] = -32'sd9925;
input_real_arr[23] = 32'sd1727;
input_real_arr[151] = 32'sd9273;
input_real_arr[87] = -32'sd7976;
input_real_arr[215] = -32'sd7997;
input_real_arr[55] = 32'sd11345;
input_real_arr[183] = 32'sd8186;
input_real_arr[119] = -32'sd10326;
input_real_arr[247] = -32'sd9488;
input_real_arr[15] = 32'sd7089;
input_real_arr[143] = 32'sd9500;
input_real_arr[79] = -32'sd6167;
input_real_arr[207] = -32'sd7846;
input_real_arr[47] = 32'sd9141;
input_real_arr[175] = 32'sd5655;
input_real_arr[111] = -32'sd13024;
input_real_arr[239] = -32'sd3910;
input_real_arr[31] = 32'sd15929;
input_real_arr[159] = 32'sd2729;
input_real_arr[95] = -32'sd19510;
input_real_arr[223] = -32'sd1595;
input_real_arr[63] = 32'sd26021;
input_real_arr[191] = 32'sd609;
input_real_arr[127] = -32'sd32767;
input_real_arr[255] = 32'sd0;
