correct_real[0] = 32'sd0; correct_imag[0] = 32'h0;
correct_real[1] = 32'sd5; correct_imag[1] = -32'h432;
correct_real[2] = 32'sd21; correct_imag[2] = -32'h868;
correct_real[3] = 32'sd47; correct_imag[3] = -32'h1301;
correct_real[4] = 32'sd85; correct_imag[4] = -32'h1730;
correct_real[5] = 32'sd134; correct_imag[5] = -32'h2188;
correct_real[6] = 32'sd193; correct_imag[6] = -32'h2617;
correct_real[7] = 32'sd264; correct_imag[7] = -32'h3069;
correct_real[8] = 32'sd344; correct_imag[8] = -32'h3499;
correct_real[9] = 32'sd440; correct_imag[9] = -32'h3970;
correct_real[10] = 32'sd547; correct_imag[10] = -32'h4436;
correct_real[11] = 32'sd667; correct_imag[11] = -32'h4916;
correct_real[12] = 32'sd800; correct_imag[12] = -32'h5399;
correct_real[13] = 32'sd950; correct_imag[13] = -32'h5906;
correct_real[14] = 32'sd1116; correct_imag[14] = -32'h6432;
correct_real[15] = 32'sd1300; correct_imag[15] = -32'h6984;
correct_real[16] = 32'sd1515; correct_imag[16] = -32'h7618;
correct_real[17] = 32'sd2186; correct_imag[17] = -32'h10329;
correct_real[18] = 32'sd2499; correct_imag[18] = -32'h11129;
correct_real[19] = 32'sd2103; correct_imag[19] = -32'h8856;
correct_real[20] = 32'sd2423; correct_imag[20] = -32'h9675;
correct_real[21] = 32'sd2787; correct_imag[21] = -32'h10577;
correct_real[22] = 32'sd4659; correct_imag[22] = -32'h16837;
correct_real[23] = 32'sd3166; correct_imag[23] = -32'h10917;
correct_real[24] = 32'sd3631; correct_imag[24] = -32'h11971;
correct_real[25] = 32'sd4078; correct_imag[25] = -32'h12873;
correct_real[26] = 32'sd4556; correct_imag[26] = -32'h13793;
correct_real[27] = 32'sd5090; correct_imag[27] = -32'h14796;
correct_real[28] = 32'sd5706; correct_imag[28] = -32'h15948;
correct_real[29] = 32'sd6468; correct_imag[29] = -32'h17402;
correct_real[30] = 32'sd7609; correct_imag[30] = -32'h19726;
correct_real[31] = 32'sd16532; correct_imag[31] = -32'h41341;
correct_real[32] = 32'sd7121; correct_imag[32] = -32'h17193;
correct_real[33] = 32'sd9100; correct_imag[33] = -32'h21229;
correct_real[34] = 32'sd11551; correct_imag[34] = -32'h26059;
correct_real[35] = 32'sd28465; correct_imag[35] = -32'h62146;
correct_real[36] = 32'sd28068; correct_imag[36] = -32'h59345;
correct_real[37] = 32'sd27248; correct_imag[37] = -32'h55828;
correct_real[38] = 32'sd5042; correct_imag[38] = -32'h10017;
correct_real[39] = 32'sd8838; correct_imag[39] = -32'h17034;
correct_real[40] = 32'sd11039; correct_imag[40] = -32'h20653;
correct_real[41] = 32'sd12946; correct_imag[41] = -32'h23522;
correct_real[42] = 32'sd14858; correct_imag[42] = -32'h26229;
correct_real[43] = 32'sd16932; correct_imag[43] = -32'h29051;
correct_real[44] = 32'sd19279; correct_imag[44] = -32'h32165;
correct_real[45] = 32'sd22070; correct_imag[45] = -32'h35818;
correct_real[46] = 32'sd25536; correct_imag[46] = -32'h40326;
correct_real[47] = 32'sd30178; correct_imag[47] = -32'h46387;
correct_real[48] = 32'sd37153; correct_imag[48] = -32'h55603;
correct_real[49] = 32'sd50679; correct_imag[49] = -32'h73867;
correct_real[50] = 32'sd140874; correct_imag[50] = -32'h200026;
correct_real[51] = 32'sd121963; correct_imag[51] = -32'h168738;
correct_real[52] = 32'sd103431; correct_imag[52] = -32'h139460;
correct_real[53] = -32'sd14053; correct_imag[53] = 32'h18470;
correct_real[54] = 32'sd12500; correct_imag[54] = -32'h16017;
correct_real[55] = 32'sd26458; correct_imag[55] = -32'h33058;
correct_real[56] = 32'sd39510; correct_imag[56] = -32'h48144;
correct_real[57] = 32'sd56304; correct_imag[57] = -32'h66915;
correct_real[58] = 32'sd87095; correct_imag[58] = -32'h100968;
correct_real[59] = 32'sd275782; correct_imag[59] = -32'h311886;
correct_real[60] = 32'sd200339; correct_imag[60] = -32'h221041;
correct_real[61] = -32'sd35281; correct_imag[61] = 32'h37979;
correct_real[62] = 32'sd30878; correct_imag[62] = -32'h32432;
correct_real[63] = 32'sd77720; correct_imag[63] = -32'h79651;
correct_real[64] = 32'sd155961; correct_imag[64] = -32'h155961;
correct_real[65] = 32'sd644199; correct_imag[65] = -32'h628579;
correct_real[66] = 32'sd165440; correct_imag[66] = -32'h157512;
correct_real[67] = 32'sd322955; correct_imag[67] = -32'h300009;
correct_real[68] = -32'sd239484; correct_imag[68] = 32'h217056;
correct_real[69] = 32'sd64157; correct_imag[69] = -32'h56730;
correct_real[70] = -32'sd190789; correct_imag[70] = 32'h164576;
correct_real[71] = -32'sd118777; correct_imag[71] = 32'h99942;
correct_real[72] = -32'sd88324; correct_imag[72] = 32'h72485;
correct_real[73] = -32'sd66722; correct_imag[73] = 32'h53401;
correct_real[74] = -32'sd45071; correct_imag[74] = 32'h35174;
correct_real[75] = -32'sd9596; correct_imag[75] = 32'h7301;
correct_real[76] = 32'sd208622; correct_imag[76] = -32'h154724;
correct_real[77] = -32'sd178346; correct_imag[77] = 32'h128908;
correct_real[78] = -32'sd105483; correct_imag[78] = 32'h74289;
correct_real[79] = -32'sd84032; correct_imag[79] = 32'h57652;
correct_real[80] = -32'sd72648; correct_imag[80] = 32'h48542;
correct_real[81] = -32'sd65024; correct_imag[81] = 32'h42303;
correct_real[82] = -32'sd59236; correct_imag[82] = 32'h37510;
correct_real[83] = -32'sd54403; correct_imag[83] = 32'h33522;
correct_real[84] = -32'sd50006; correct_imag[84] = 32'h29972;
correct_real[85] = -32'sd45547; correct_imag[85] = 32'h26545;
correct_real[86] = -32'sd40204; correct_imag[86] = 32'h22775;
correct_real[87] = -32'sd31440; correct_imag[87] = 32'h17304;
correct_real[88] = 32'sd9862; correct_imag[88] = -32'h5271;
correct_real[89] = -32'sd59793; correct_imag[89] = 32'h31023;
correct_real[90] = -32'sd10724; correct_imag[90] = 32'h5398;
correct_real[91] = -32'sd65117; correct_imag[91] = 32'h31782;
correct_real[92] = -32'sd24384; correct_imag[92] = 32'h11532;
correct_real[93] = -32'sd70699; correct_imag[93] = 32'h32382;
correct_real[94] = -32'sd56213; correct_imag[94] = 32'h24917;
correct_real[95] = -32'sd51204; correct_imag[95] = 32'h21949;
correct_real[96] = -32'sd48155; correct_imag[96] = 32'h19946;
correct_real[97] = -32'sd45809; correct_imag[97] = 32'h18319;
correct_real[98] = -32'sd43675; correct_imag[98] = 32'h16847;
correct_real[99] = -32'sd40988; correct_imag[99] = 32'h15236;
correct_real[100] = -32'sd31257; correct_imag[100] = 32'h11184;
correct_real[101] = -32'sd50156; correct_imag[101] = 32'h17254;
correct_real[102] = -32'sd44516; correct_imag[102] = 32'h14706;
correct_real[103] = -32'sd42667; correct_imag[103] = 32'h13517;
correct_real[104] = -32'sd41516; correct_imag[104] = 32'h12593;
correct_real[105] = -32'sd40633; correct_imag[105] = 32'h11783;
correct_real[106] = -32'sd39910; correct_imag[106] = 32'h11044;
correct_real[107] = -32'sd39276; correct_imag[107] = 32'h10352;
correct_real[108] = -32'sd38670; correct_imag[108] = 32'h9686;
correct_real[109] = -32'sd38087; correct_imag[109] = 32'h9045;
correct_real[110] = -32'sd37394; correct_imag[110] = 32'h8397;
correct_real[111] = -32'sd35712; correct_imag[111] = 32'h7560;
correct_real[112] = -32'sd37219; correct_imag[112] = 32'h7403;
correct_real[113] = -32'sd37694; correct_imag[113] = 32'h7018;
correct_real[114] = -32'sd38352; correct_imag[114] = 32'h6654;
correct_real[115] = -32'sd37399; correct_imag[115] = 32'h6017;
correct_real[116] = -32'sd36970; correct_imag[116] = 32'h5484;
correct_real[117] = -32'sd36644; correct_imag[117] = 32'h4976;
correct_real[118] = -32'sd36292; correct_imag[118] = 32'h4476;
correct_real[119] = -32'sd36424; correct_imag[119] = 32'h4039;
correct_real[120] = -32'sd36164; correct_imag[120] = 32'h3561;
correct_real[121] = -32'sd36000; correct_imag[121] = 32'h3100;
correct_real[122] = -32'sd35872; correct_imag[122] = 32'h2646;
correct_real[123] = -32'sd35764; correct_imag[123] = 32'h2197;
correct_real[124] = -32'sd35678; correct_imag[124] = 32'h1752;
correct_real[125] = -32'sd35641; correct_imag[125] = 32'h1312;
correct_real[126] = -32'sd35595; correct_imag[126] = 32'h873;
correct_real[127] = -32'sd35568; correct_imag[127] = 32'h436;
correct_real[128] = -32'sd35550; correct_imag[128] = 32'h0;
correct_real[129] = -32'sd35568; correct_imag[129] = -32'h436;
correct_real[130] = -32'sd35595; correct_imag[130] = -32'h873;
correct_real[131] = -32'sd35641; correct_imag[131] = -32'h1312;
correct_real[132] = -32'sd35678; correct_imag[132] = -32'h1752;
correct_real[133] = -32'sd35764; correct_imag[133] = -32'h2197;
correct_real[134] = -32'sd35872; correct_imag[134] = -32'h2646;
correct_real[135] = -32'sd36000; correct_imag[135] = -32'h3100;
correct_real[136] = -32'sd36164; correct_imag[136] = -32'h3561;
correct_real[137] = -32'sd36424; correct_imag[137] = -32'h4039;
correct_real[138] = -32'sd36292; correct_imag[138] = -32'h4476;
correct_real[139] = -32'sd36644; correct_imag[139] = -32'h4976;
correct_real[140] = -32'sd36970; correct_imag[140] = -32'h5484;
correct_real[141] = -32'sd37399; correct_imag[141] = -32'h6017;
correct_real[142] = -32'sd38352; correct_imag[142] = -32'h6654;
correct_real[143] = -32'sd37694; correct_imag[143] = -32'h7018;
correct_real[144] = -32'sd37219; correct_imag[144] = -32'h7403;
correct_real[145] = -32'sd35712; correct_imag[145] = -32'h7560;
correct_real[146] = -32'sd37394; correct_imag[146] = -32'h8397;
correct_real[147] = -32'sd38087; correct_imag[147] = -32'h9045;
correct_real[148] = -32'sd38670; correct_imag[148] = -32'h9686;
correct_real[149] = -32'sd39276; correct_imag[149] = -32'h10352;
correct_real[150] = -32'sd39910; correct_imag[150] = -32'h11044;
correct_real[151] = -32'sd40633; correct_imag[151] = -32'h11783;
correct_real[152] = -32'sd41516; correct_imag[152] = -32'h12593;
correct_real[153] = -32'sd42667; correct_imag[153] = -32'h13517;
correct_real[154] = -32'sd44516; correct_imag[154] = -32'h14706;
correct_real[155] = -32'sd50156; correct_imag[155] = -32'h17254;
correct_real[156] = -32'sd31257; correct_imag[156] = -32'h11184;
correct_real[157] = -32'sd40988; correct_imag[157] = -32'h15236;
correct_real[158] = -32'sd43675; correct_imag[158] = -32'h16847;
correct_real[159] = -32'sd45809; correct_imag[159] = -32'h18319;
correct_real[160] = -32'sd48155; correct_imag[160] = -32'h19946;
correct_real[161] = -32'sd51204; correct_imag[161] = -32'h21949;
correct_real[162] = -32'sd56213; correct_imag[162] = -32'h24917;
correct_real[163] = -32'sd70699; correct_imag[163] = -32'h32382;
correct_real[164] = -32'sd24384; correct_imag[164] = -32'h11532;
correct_real[165] = -32'sd65117; correct_imag[165] = -32'h31782;
correct_real[166] = -32'sd10724; correct_imag[166] = -32'h5398;
correct_real[167] = -32'sd59793; correct_imag[167] = -32'h31023;
correct_real[168] = 32'sd9862; correct_imag[168] = 32'h5271;
correct_real[169] = -32'sd31440; correct_imag[169] = -32'h17304;
correct_real[170] = -32'sd40204; correct_imag[170] = -32'h22775;
correct_real[171] = -32'sd45547; correct_imag[171] = -32'h26545;
correct_real[172] = -32'sd50006; correct_imag[172] = -32'h29972;
correct_real[173] = -32'sd54403; correct_imag[173] = -32'h33522;
correct_real[174] = -32'sd59236; correct_imag[174] = -32'h37510;
correct_real[175] = -32'sd65024; correct_imag[175] = -32'h42303;
correct_real[176] = -32'sd72648; correct_imag[176] = -32'h48542;
correct_real[177] = -32'sd84032; correct_imag[177] = -32'h57652;
correct_real[178] = -32'sd105483; correct_imag[178] = -32'h74289;
correct_real[179] = -32'sd178346; correct_imag[179] = -32'h128908;
correct_real[180] = 32'sd208622; correct_imag[180] = 32'h154724;
correct_real[181] = -32'sd9596; correct_imag[181] = -32'h7301;
correct_real[182] = -32'sd45071; correct_imag[182] = -32'h35174;
correct_real[183] = -32'sd66722; correct_imag[183] = -32'h53401;
correct_real[184] = -32'sd88324; correct_imag[184] = -32'h72485;
correct_real[185] = -32'sd118777; correct_imag[185] = -32'h99942;
correct_real[186] = -32'sd190789; correct_imag[186] = -32'h164576;
correct_real[187] = 32'sd64157; correct_imag[187] = 32'h56730;
correct_real[188] = -32'sd239484; correct_imag[188] = -32'h217056;
correct_real[189] = 32'sd322955; correct_imag[189] = 32'h300009;
correct_real[190] = 32'sd165440; correct_imag[190] = 32'h157512;
correct_real[191] = 32'sd644199; correct_imag[191] = 32'h628579;
correct_real[192] = 32'sd155961; correct_imag[192] = 32'h155961;
correct_real[193] = 32'sd77720; correct_imag[193] = 32'h79651;
correct_real[194] = 32'sd30878; correct_imag[194] = 32'h32432;
correct_real[195] = -32'sd35281; correct_imag[195] = -32'h37979;
correct_real[196] = 32'sd200339; correct_imag[196] = 32'h221041;
correct_real[197] = 32'sd275782; correct_imag[197] = 32'h311886;
correct_real[198] = 32'sd87095; correct_imag[198] = 32'h100968;
correct_real[199] = 32'sd56304; correct_imag[199] = 32'h66915;
correct_real[200] = 32'sd39510; correct_imag[200] = 32'h48144;
correct_real[201] = 32'sd26458; correct_imag[201] = 32'h33058;
correct_real[202] = 32'sd12500; correct_imag[202] = 32'h16017;
correct_real[203] = -32'sd14053; correct_imag[203] = -32'h18470;
correct_real[204] = 32'sd103431; correct_imag[204] = 32'h139460;
correct_real[205] = 32'sd121963; correct_imag[205] = 32'h168738;
correct_real[206] = 32'sd140874; correct_imag[206] = 32'h200026;
correct_real[207] = 32'sd50679; correct_imag[207] = 32'h73867;
correct_real[208] = 32'sd37153; correct_imag[208] = 32'h55603;
correct_real[209] = 32'sd30178; correct_imag[209] = 32'h46387;
correct_real[210] = 32'sd25536; correct_imag[210] = 32'h40326;
correct_real[211] = 32'sd22070; correct_imag[211] = 32'h35818;
correct_real[212] = 32'sd19279; correct_imag[212] = 32'h32165;
correct_real[213] = 32'sd16932; correct_imag[213] = 32'h29051;
correct_real[214] = 32'sd14858; correct_imag[214] = 32'h26229;
correct_real[215] = 32'sd12946; correct_imag[215] = 32'h23522;
correct_real[216] = 32'sd11039; correct_imag[216] = 32'h20653;
correct_real[217] = 32'sd8838; correct_imag[217] = 32'h17034;
correct_real[218] = 32'sd5042; correct_imag[218] = 32'h10017;
correct_real[219] = 32'sd27248; correct_imag[219] = 32'h55828;
correct_real[220] = 32'sd28068; correct_imag[220] = 32'h59345;
correct_real[221] = 32'sd28465; correct_imag[221] = 32'h62146;
correct_real[222] = 32'sd11551; correct_imag[222] = 32'h26059;
correct_real[223] = 32'sd9100; correct_imag[223] = 32'h21229;
correct_real[224] = 32'sd7121; correct_imag[224] = 32'h17193;
correct_real[225] = 32'sd16532; correct_imag[225] = 32'h41341;
correct_real[226] = 32'sd7609; correct_imag[226] = 32'h19726;
correct_real[227] = 32'sd6468; correct_imag[227] = 32'h17402;
correct_real[228] = 32'sd5706; correct_imag[228] = 32'h15948;
correct_real[229] = 32'sd5090; correct_imag[229] = 32'h14796;
correct_real[230] = 32'sd4556; correct_imag[230] = 32'h13793;
correct_real[231] = 32'sd4078; correct_imag[231] = 32'h12873;
correct_real[232] = 32'sd3631; correct_imag[232] = 32'h11971;
correct_real[233] = 32'sd3166; correct_imag[233] = 32'h10917;
correct_real[234] = 32'sd4659; correct_imag[234] = 32'h16837;
correct_real[235] = 32'sd2787; correct_imag[235] = 32'h10577;
correct_real[236] = 32'sd2423; correct_imag[236] = 32'h9675;
correct_real[237] = 32'sd2103; correct_imag[237] = 32'h8856;
correct_real[238] = 32'sd2499; correct_imag[238] = 32'h11129;
correct_real[239] = 32'sd2186; correct_imag[239] = 32'h10329;
correct_real[240] = 32'sd1515; correct_imag[240] = 32'h7618;
correct_real[241] = 32'sd1300; correct_imag[241] = 32'h6984;
correct_real[242] = 32'sd1116; correct_imag[242] = 32'h6432;
correct_real[243] = 32'sd950; correct_imag[243] = 32'h5906;
correct_real[244] = 32'sd800; correct_imag[244] = 32'h5399;
correct_real[245] = 32'sd667; correct_imag[245] = 32'h4916;
correct_real[246] = 32'sd547; correct_imag[246] = 32'h4436;
correct_real[247] = 32'sd440; correct_imag[247] = 32'h3970;
correct_real[248] = 32'sd344; correct_imag[248] = 32'h3499;
correct_real[249] = 32'sd264; correct_imag[249] = 32'h3069;
correct_real[250] = 32'sd193; correct_imag[250] = 32'h2617;
correct_real[251] = 32'sd134; correct_imag[251] = 32'h2188;
correct_real[252] = 32'sd85; correct_imag[252] = 32'h1730;
correct_real[253] = 32'sd47; correct_imag[253] = 32'h1301;
correct_real[254] = 32'sd21; correct_imag[254] = 32'h868;
correct_real[255] = 32'sd5; correct_imag[255] = 32'h432;
