correct_real[0] = 32'sd0; correct_imag[0] = 32'h0;
correct_real[1] = 32'sd77; correct_imag[1] = -32'h1584;
correct_real[2] = 32'sd320; correct_imag[2] = -32'h3253;
correct_real[3] = 32'sd821; correct_imag[3] = -32'h5536;
correct_real[4] = 32'sd1594; correct_imag[4] = -32'h8014;
correct_real[5] = 32'sd3233; correct_imag[5] = -32'h12909;
correct_real[6] = 32'sd3009; correct_imag[6] = -32'h9920;
correct_real[7] = 32'sd4506; correct_imag[7] = -32'h12594;
correct_real[8] = 32'sd6469; correct_imag[8] = -32'h15618;
correct_real[9] = 32'sd9211; correct_imag[9] = -32'h19476;
correct_real[10] = 32'sd13361; correct_imag[10] = -32'h24998;
correct_real[11] = 32'sd21172; correct_imag[11] = -32'h35324;
correct_real[12] = 32'sd75161; correct_imag[12] = -32'h112486;
correct_real[13] = 32'sd11937; correct_imag[13] = -32'h16095;
correct_real[14] = 32'sd36224; correct_imag[14] = -32'h44139;
correct_real[15] = 32'sd125355; correct_imag[15] = -32'h138308;
correct_real[16] = 32'sd130035; correct_imag[16] = -32'h130035;
correct_real[17] = 32'sd152429; correct_imag[17] = -32'h138153;
correct_real[18] = 32'sd50467; correct_imag[18] = -32'h41417;
correct_real[19] = -32'sd51918; correct_imag[19] = 32'h38505;
correct_real[20] = -32'sd49736; correct_imag[20] = 32'h33233;
correct_real[21] = -32'sd73406; correct_imag[21] = 32'h43997;
correct_real[22] = -32'sd22680; correct_imag[22] = 32'h12123;
correct_real[23] = -32'sd71072; correct_imag[23] = 32'h33614;
correct_real[24] = -32'sd47509; correct_imag[24] = 32'h19679;
correct_real[25] = -32'sd53211; correct_imag[25] = 32'h19039;
correct_real[26] = -32'sd44499; correct_imag[26] = 32'h13498;
correct_real[27] = -32'sd44479; correct_imag[27] = 32'h11141;
correct_real[28] = -32'sd42454; correct_imag[28] = 32'h8444;
correct_real[29] = -32'sd42871; correct_imag[29] = 32'h6359;
correct_real[30] = -32'sd41083; correct_imag[30] = 32'h4046;
correct_real[31] = -32'sd40379; correct_imag[31] = 32'h1983;
correct_real[32] = -32'sd40174; correct_imag[32] = 32'h0;
correct_real[33] = -32'sd40379; correct_imag[33] = -32'h1983;
correct_real[34] = -32'sd41083; correct_imag[34] = -32'h4046;
correct_real[35] = -32'sd42871; correct_imag[35] = -32'h6359;
correct_real[36] = -32'sd42454; correct_imag[36] = -32'h8444;
correct_real[37] = -32'sd44479; correct_imag[37] = -32'h11141;
correct_real[38] = -32'sd44499; correct_imag[38] = -32'h13498;
correct_real[39] = -32'sd53211; correct_imag[39] = -32'h19039;
correct_real[40] = -32'sd47509; correct_imag[40] = -32'h19679;
correct_real[41] = -32'sd71072; correct_imag[41] = -32'h33614;
correct_real[42] = -32'sd22680; correct_imag[42] = -32'h12123;
correct_real[43] = -32'sd73406; correct_imag[43] = -32'h43997;
correct_real[44] = -32'sd49736; correct_imag[44] = -32'h33233;
correct_real[45] = -32'sd51918; correct_imag[45] = -32'h38505;
correct_real[46] = 32'sd50467; correct_imag[46] = 32'h41417;
correct_real[47] = 32'sd152429; correct_imag[47] = 32'h138153;
correct_real[48] = 32'sd130035; correct_imag[48] = 32'h130035;
correct_real[49] = 32'sd125355; correct_imag[49] = 32'h138308;
correct_real[50] = 32'sd36224; correct_imag[50] = 32'h44139;
correct_real[51] = 32'sd11937; correct_imag[51] = 32'h16095;
correct_real[52] = 32'sd75161; correct_imag[52] = 32'h112486;
correct_real[53] = 32'sd21172; correct_imag[53] = 32'h35324;
correct_real[54] = 32'sd13361; correct_imag[54] = 32'h24998;
correct_real[55] = 32'sd9211; correct_imag[55] = 32'h19476;
correct_real[56] = 32'sd6469; correct_imag[56] = 32'h15618;
correct_real[57] = 32'sd4506; correct_imag[57] = 32'h12594;
correct_real[58] = 32'sd3009; correct_imag[58] = 32'h9920;
correct_real[59] = 32'sd3233; correct_imag[59] = 32'h12909;
correct_real[60] = 32'sd1594; correct_imag[60] = 32'h8014;
correct_real[61] = 32'sd821; correct_imag[61] = 32'h5536;
correct_real[62] = 32'sd320; correct_imag[62] = 32'h3253;
correct_real[63] = 32'sd77; correct_imag[63] = 32'h1584;
