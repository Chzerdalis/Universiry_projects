input_real[0] = 32'sd0;
input_real[1] = 32'sd32514;
input_real[2] = -32'sd13903;
input_real[3] = -32'sd25330;
input_real[4] = 32'sd26358;
input_real[5] = 32'sd14680;
input_real[6] = -32'sd32175;
input_real[7] = -32'sd183;
input_real[8] = 32'sd31853;
input_real[9] = -32'sd14879;
input_real[10] = -32'sd26385;
input_real[11] = 32'sd25483;
input_real[12] = 32'sd14197;
input_real[13] = -32'sd32149;
input_real[14] = 32'sd346;
input_real[15] = 32'sd32758;
input_real[16] = -32'sd13820;
input_real[17] = -32'sd25429;
input_real[18] = 32'sd26102;
input_real[19] = 32'sd14329;
input_real[20] = -32'sd32536;
input_real[21] = -32'sd465;
input_real[22] = 32'sd31719;
input_real[23] = -32'sd14833;
input_real[24] = -32'sd26170;
input_real[25] = 32'sd25814;
input_real[26] = 32'sd14565;
input_real[27] = -32'sd31835;
input_real[28] = 32'sd530;
input_real[29] = 32'sd32767;
input_real[30] = -32'sd13989;
input_real[31] = -32'sd25734;
input_real[32] = 32'sd25734;
input_real[33] = 32'sd13989;
input_real[34] = -32'sd32767;
input_real[35] = -32'sd530;
input_real[36] = 32'sd31835;
input_real[37] = -32'sd14565;
input_real[38] = -32'sd25814;
input_real[39] = 32'sd26170;
input_real[40] = 32'sd14833;
input_real[41] = -32'sd31719;
input_real[42] = 32'sd465;
input_real[43] = 32'sd32536;
input_real[44] = -32'sd14329;
input_real[45] = -32'sd26102;
input_real[46] = 32'sd25429;
input_real[47] = 32'sd13820;
input_real[48] = -32'sd32758;
input_real[49] = -32'sd346;
input_real[50] = 32'sd32149;
input_real[51] = -32'sd14197;
input_real[52] = -32'sd25483;
input_real[53] = 32'sd26385;
input_real[54] = 32'sd14879;
input_real[55] = -32'sd31853;
input_real[56] = 32'sd183;
input_real[57] = 32'sd32175;
input_real[58] = -32'sd14680;
input_real[59] = -32'sd26358;
input_real[60] = 32'sd25330;
input_real[61] = 32'sd13903;
input_real[62] = -32'sd32514;
input_real[63] = 32'sd0;
